/*
     __        __   __   ___ ___ ___  __  
    |__)  /\  |__) |__) |__   |   |  /  \ 
    |    /~~\ |  \ |  \ |___  |   |  \__/ 


    Module: DP Package
    (c) 2021, 2022 by Parretto B.V.

    History
    =======
    v1.0 - Initial release

    License
    =======
    This License will apply to the use of the IP-core (as defined in the License). 
    Please read the License carefully so that you know what your rights and obligations are when using the IP-core.
    The acceptance of this License constitutes a valid and binding agreement between Parretto and you for the use of the IP-core. 
    If you download and/or make any use of the IP-core you agree to be bound by this License. 
    The License is available for download and print at www.parretto.com/license.html
    Parretto grants you, as the Licensee, a free, non-exclusive, non-transferable, limited right to use the IP-core 
    solely for internal business purposes for the term and conditions of the License. 
    You are also allowed to create Modifications for internal business purposes, but explicitly only under the conditions of art. 3.2.
    You are, however, obliged to pay the License Fees to Parretto for the use of the IP-core, or any Modification, in, or embodied in, 
    a physical or non-tangible product or service that has substantial commercial, industrial or non-consumer uses. 
*/

package prt_dp_pkg;

// Parameters

// Symbols
localparam P_SYM_BS = 'h1_bc;	// K28.5
localparam P_SYM_BF = 'h1_7c;	// K28.3
localparam P_SYM_BE = 'h1_fb;	// K27.7
localparam P_SYM_FS = 'h1_fe;	// K30.7
localparam P_SYM_FE = 'h1_f7;	// K23.7
localparam P_SYM_SR = 'h1_1c;	// K28.0
localparam P_SYM_SS = 'h1_5c;	// K28.2
localparam P_SYM_SE = 'h1_fd;	// K29.7

endpackage
